// Copyright (c) 2015 Cornell University.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

/* DO NOT MODIFY, AUTO GENERATED BY P4 COMPILER */

import BuildVector::*;
import DefaultValue::*;
import FIFOF::*;
import GetPut::*;
import Pipe::*;
import StmtFSM::*;
import SpecialFIFOs::*;
import Vector::*;

import Ethernet::*;
import Types::*;

interface Parser;
   method Action enqPacketData(EtherData b);
   method Action parserReset();
   interface PipeOut#(void) parseDone;
   interface PipeOut#(PHV_port_mapping) phvOut;
   interface PipeOut#(Bit#(128)) payloadOut;
endinterface

(* synthesize *)
module mkParser(Parser);

   Reg#(Bit#(32)) cycle <- mkReg(0);
   FIFOF#(EtherData) data_fifo_in <- mkSizedFIFOF(1);
   FIFOF#(Bit#(128)) header_fifo_in <- mkSizedFIFOF(1);
   FIFOF#(Bit#(16)) parse_ethernet_fifo_out <- mkSizedFIFOF(1);
   FIFOF#(Bit#(144)) parse_ipv4_fifo_0 <- mkSizedFIFOF(1);
   FIFOF#(Bit#(112)) parse_ipv4_fifo_out <- mkSizedFIFOF(1);
   FIFOF#(void) parse_done_fifo <- mkSizedFIFOF(1);
   FIFOF#(void) payload_cfFifo <- mkSizedFIFOF(1);

   Reg#(HeaderType_ethernet) reg_ethernet <- mkReg(defaultValue);
   Reg#(HeaderType_ipv4) reg_ipv4 <- mkReg(defaultValue);
   Reg#(HeaderType_standard_metadata) reg_standard_metadata <- mkReg(defaultValue);
   Reg#(HeaderType_ingress_metadata) reg_ingress_metadata <- mkReg(defaultValue);

   FIFOF#(PHV_port_mapping) fifo_out_phv <- mkBypassFIFOF();
   FIFOF#(Bit#(128)) fifo_out_payload <- mkBypassFIFOF();

   rule every;
      cycle <= cycle + 1;
   endrule

   // One Stmt that says it all
   Stmt parseSeq =
   seq
   action // parse_ethernet
      let data <- toGet(header_fifo_in).get;
      Vector#(128, Bit#(1)) dataVec = unpack(data);
      Vector#(48, Bit#(1)) dstAddr = takeAt(0, dataVec);
      Vector#(48, Bit#(1)) srcAddr = takeAt(48, dataVec);
      Vector#(16, Bit#(1)) etherType = takeAt(96, dataVec);
      Vector#(16, Bit#(1)) residue = takeAt(112, dataVec);
      HeaderType_ethernet ethernet = defaultValue;
      ethernet.dstAddr = pack(dstAddr);
      ethernet.srcAddr = pack(srcAddr);
      ethernet.etherType = pack(etherType);
      reg_ethernet <= ethernet;
      parse_ethernet_fifo_out.enq(pack(residue));
      $display("parse ethernet");
   endaction
   action // parse_ipv4
      let data_current <- toGet(header_fifo_in).get;
      let residue_last <- toGet(parse_ethernet_fifo_out).get;
      Bit#(144) data = {data_current, residue_last};
      Vector#(144, Bit#(1)) dataVec = unpack(data);
      parse_ipv4_fifo_0.enq(data);
      $display("wait for ip");
   endaction
   action // parse_ipv4 0
      let data_current <- toGet(header_fifo_in).get;
      let data_delayed <- toGet(parse_ipv4_fifo_0).get;
      Bit#(272) data = {data_current, data_delayed};
      Vector#(272, Bit#(1)) dataVec = unpack(data);
      Vector#(4, Bit#(1)) version = takeAt(0, dataVec);
      Vector#(4, Bit#(1)) ihl = takeAt(4, dataVec);
      Vector#(8, Bit#(1)) diffserv = takeAt(8, dataVec);
      Vector#(16, Bit#(1)) totalLen = takeAt(16, dataVec);
      Vector#(16, Bit#(1)) identification = takeAt(32, dataVec);
      Vector#(3, Bit#(1)) flags = takeAt(48, dataVec);
      Vector#(13, Bit#(1)) fragOffset = takeAt(51, dataVec);
      Vector#(8, Bit#(1)) ttl = takeAt(64, dataVec);
      Vector#(8, Bit#(1)) protocol = takeAt(72, dataVec);
      Vector#(16, Bit#(1)) hdrChecksum = takeAt(80, dataVec);
      Vector#(32, Bit#(1)) srcAddr = takeAt(96, dataVec);
      Vector#(32, Bit#(1)) dstAddr = takeAt(128, dataVec);
      Vector#(112, Bit#(1)) residue = takeAt(160, dataVec);
      HeaderType_ipv4 ipv4 = defaultValue;
      ipv4.version = pack(version);
      ipv4.ihl = pack(ihl);
      ipv4.diffserv = pack(diffserv);
      ipv4.totalLen = pack(totalLen);
      ipv4.identification = pack(identification);
      ipv4.flags = pack(flags);
      ipv4.fragOffset = pack(fragOffset);
      ipv4.ttl = pack(ttl);
      ipv4.protocol = pack(protocol);
      ipv4.hdrChecksum = pack(hdrChecksum);
      ipv4.srcAddr = pack(srcAddr);
      ipv4.dstAddr = pack(dstAddr);
      reg_ipv4 <= ipv4;
      parse_done_fifo.enq(?);

      PHV_port_mapping phv = defaultValue;
      phv.ipv4_dstAddr = ipv4.dstAddr;
      fifo_out_phv.enq(phv);
      payload_cfFifo.enq(?);
   endaction
   endseq;

   // control parsing FSM
   FSM parseFSM <- mkFSM(parseSeq);
   Once parseOnce <- mkOnce(parseFSM.start);

   rule parse_starts;
      parseOnce.start;
   endrule

   rule forward_header (!payload_cfFifo.notEmpty);
      let v <- toGet(data_fifo_in).get;
      header_fifo_in.enq(v.data);
      fifo_out_payload.enq(v.data);
   endrule

   rule forward_payload (payload_cfFifo.notEmpty);
      let v <- toGet(data_fifo_in).get;
      fifo_out_payload.enq(v.data);
      if (v.eop) begin
         payload_cfFifo.deq;
      end
   endrule

   method Action parserReset();
      parseOnce.clear;
   endmethod

   method Action enqPacketData(EtherData b);
      $display("enqueue packet data %x", b);
      data_fifo_in.enq(b);
   endmethod

   interface parseDone = toPipeOut(parse_done_fifo);
   interface phvOut = toPipeOut(fifo_out_phv);
   interface payloadOut = toPipeOut(fifo_out_payload);
endmodule

