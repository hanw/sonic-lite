// Copyright (c) 2015 Cornell University.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

/* DO NOT MODIFY, AUTO GENERATED BY P4 COMPILER */

import BuildVector::*;
import Connectable::*;
import DefaultValue::*;
import FIFO::*;
import FIFOF::*;
import FShow::*;
import GetPut::*;
import Pipe::*;
import StmtFSM::*;
import SpecialFIFOs::*;
import Vector::*;

import Ethernet::*;
import Types::*;

interface Parser;
   // derive parseReset from start of packet
   method Action parserReset();
   interface PipeIn#(EtherData) frameIn;
   interface PipeOut#(void) parseDone;
   interface PipeOut#(PHV_port_mapping) phvOut;
   interface PipeOut#(Bit#(128)) payloadOut;
endinterface

interface ParseEthernet;
   interface PipeIn#(Bit#(128)) packetIn;
   interface PipeOut#(Ethernet_t) parsedOut;
   interface PipeOut#(Bit#(16)) unparsedOut; // number is parse state id
   interface PipeOut#(Bit#(16)) nextState; // upon completion, tell where to send new data.
   interface PipeIn#(Bool) start;
   interface PipeOut#(Bool) done;
   method Action init;
   method Action clear;
endinterface

interface ParseVlan;
   interface PipeIn#(Bit#(128)) packetIn;
   interface PipeOut#(Vlan_tag_t) parsedOut;
   interface PipeOut#(Bit#(16)) unparsedOut;
   interface PipeIn#(Bool) start;
   interface PipeOut#(Bool) done;
   method Action init;
   method Action clear;
endinterface

interface ParseIpv4;
   interface PipeIn#(Bit#(128)) packetIn;
   interface PipeIn#(Bit#(16)) unparsedIn;
   interface PipeOut#(Ipv4_t) parsedOut;
   interface PipeOut#(Bit#(112)) unparsedOut;
   interface PipeOut#(Bit#(16)) nextState; // upon completion, tell where to send new data.
   interface PipeIn#(Bool) start;
   interface PipeOut#(Bool) done;
   method Action init;
   method Action clear;
endinterface

module mkParseEthernet(ParseEthernet);
   FIFOF#(Bool) start_fifo <- mkBypassFIFOF;
   FIFOF#(Bit#(128)) packet_in_fifo <- mkBypassFIFOF;
   FIFOF#(Ethernet_t) parsed_out_fifo <- mkSizedFIFOF(1);
   FIFOF#(Bit#(16))  unparsed_out_fifo <- mkSizedFIFOF(1);
   FIFOF#(Bool) finish_fifo <- mkBypassFIFOF;

   let verbose = True;
   Reg#(Cycle_t) cycle <- mkReg(0);
   rule every;
      cycle <= cycle + 1;
   endrule

   Stmt parse_ethernet =
   seq
   action // parse_ethernet
      let data <- toGet(packet_in_fifo).get;
      Vector#(128, Bit#(1)) dataVec = unpack(data);
      Vector#(48, Bit#(1)) dstAddr = takeAt(0, dataVec);
      Vector#(48, Bit#(1)) srcAddr = takeAt(48, dataVec);
      Vector#(16, Bit#(1)) etherType = takeAt(96, dataVec);
      Vector#(16, Bit#(1)) unparsed = takeAt(112, dataVec);
      Ethernet_t ethernet = defaultValue;
      ethernet.dstAddr = pack(dstAddr);
      ethernet.srcAddr = pack(srcAddr);
      ethernet.etherType = pack(etherType);
      if (verbose) $display(fshow(cycle)
                            +fshow("ether.dstAddr=")+fshow(ethernet.dstAddr)
                            +fshow("ether.srcAddr=")+fshow(ethernet.srcAddr));
      finish_fifo.enq(True);
   endaction
   endseq;

   FSM fsm_parse_ethernet <- mkFSMWithPred(parse_ethernet, True);
   Once once_parse_ethernet <- mkOnce(fsm_parse_ethernet.start);

   method Action init = once_parse_ethernet.start;
   method Action clear = once_parse_ethernet.clear;
   interface done = toPipeOut(finish_fifo);
   interface packetIn = toPipeIn(packet_in_fifo);
   interface unparsedOut = toPipeOut(unparsed_out_fifo);
   interface parsedOut = toPipeOut(parsed_out_fifo);
   interface start = toPipeIn(start_fifo);
endmodule

module mkParseVlan(ParseVlan);
   FIFOF#(Bool) start_fifo <- mkBypassFIFOF;
   FIFOF#(Bit#(128)) packet_in_fifo <- mkBypassFIFOF;
   FIFOF#(Vlan_tag_t) parsed_out_fifo <- mkSizedFIFOF(1);
   FIFOF#(Bit#(16)) unparsed_out_fifo <- mkSizedFIFOF(1);
   FIFOF#(Bool) finish_fifo <- mkBypassFIFOF;

   let verbose = True;
   Reg#(Cycle_t) cycle <- mkReg(0);
   rule every;
      cycle <= cycle + 1;
   endrule

   Stmt parse_vlan =
   seq
   action
   noAction;
   endaction
   endseq;

endmodule

module mkParseIpv4(ParseIpv4);
   FIFOF#(Bool) start_fifo <- mkBypassFIFOF;
   FIFOF#(Bool) done_fifo <- mkBypassFIFOF;
   FIFOF#(Bit#(128)) packet_in_fifo <- mkBypassFIFOF;
   FIFOF#(Ipv4_t) parsed_out_fifo <- mkSizedFIFOF(1);
   FIFOF#(Bit#(16)) unparsed_in_fifo <- mkBypassFIFOF;
   FIFOF#(Bit#(112)) unparsed_out_fifo <- mkSizedFIFOF(1);
   FIFOF#(Bit#(144)) internal_fifo <- mkSizedFIFOF(1);

   let verbose = True;
   Reg#(Cycle_t) cycle <- mkReg(0);
   rule every;
      cycle <= cycle + 1;
   endrule

   // Can we use List#() to simplify design??
   // We need a collection for fields to extract. not all fields are required.
   Stmt parse_ipv4 =
   seq
   action // parse_ipv4
      let data_current <- toGet(packet_in_fifo).get;
      //let residue_last <- toGet(unparsed_in_fifo).get;
      Bit#(144) data = {data_current, 0}; //residue_last};
      Vector#(144, Bit#(1)) dataVec = unpack(data);
      internal_fifo.enq(data);
      if (verbose) $display(fshow(cycle) + fshow("wait one cycle!"));
   endaction
   action // parse_ipv4 0
      let data_current <- toGet(packet_in_fifo).get;
      let data_delayed <- toGet(internal_fifo).get;
      Bit#(272) data = {data_current, data_delayed};
      Vector#(272, Bit#(1)) dataVec = unpack(data);
      Vector#(4, Bit#(1)) version = takeAt(0, dataVec);
      Vector#(4, Bit#(1)) ihl = takeAt(4, dataVec);
      Vector#(8, Bit#(1)) diffserv = takeAt(8, dataVec);
      Vector#(16, Bit#(1)) totalLen = takeAt(16, dataVec);
      Vector#(16, Bit#(1)) identification = takeAt(32, dataVec);
      Vector#(3, Bit#(1)) flags = takeAt(48, dataVec);
      Vector#(13, Bit#(1)) fragOffset = takeAt(51, dataVec);
      Vector#(8, Bit#(1)) ttl = takeAt(64, dataVec);
      Vector#(8, Bit#(1)) protocol = takeAt(72, dataVec);
      Vector#(16, Bit#(1)) hdrChecksum = takeAt(80, dataVec);
      Vector#(32, Bit#(1)) srcAddr = takeAt(96, dataVec);
      Vector#(32, Bit#(1)) dstAddr = takeAt(128, dataVec);
      Vector#(112, Bit#(1)) residue = takeAt(160, dataVec);
      Ipv4_t ipv4 = defaultValue;
      ipv4.version = pack(version);
      ipv4.ihl = pack(ihl);
      ipv4.diffserv = pack(diffserv);
      ipv4.totalLen = pack(totalLen);
      ipv4.identification = pack(identification);
      ipv4.flags = pack(flags);
      ipv4.fragOffset = pack(fragOffset);
      ipv4.ttl = pack(ttl);
      ipv4.protocol = pack(protocol);
      ipv4.hdrChecksum = pack(hdrChecksum);
      ipv4.srcAddr = pack(srcAddr);
      ipv4.dstAddr = pack(dstAddr);
      if (verbose) $display(fshow(cycle)
                            +fshow("ipv4.dstAddr=")+fshow(ipv4.dstAddr)
                            +fshow("ipv4.srcAddr=")+fshow(ipv4.srcAddr));
      done_fifo.enq(True);
   endaction
   endseq;

   FSM fsm_parse_ipv4 <- mkFSMWithPred(parse_ipv4, True);
   Once once_parse_ipv4 <- mkOnce(fsm_parse_ipv4.start);

   method Action init = once_parse_ipv4.start;
   method Action clear = once_parse_ipv4.clear;
   interface packetIn = toPipeIn(packet_in_fifo);
   interface unparsedIn = toPipeIn(unparsed_in_fifo);
   interface unparsedOut = toPipeOut(unparsed_out_fifo);
   interface parsedOut = toPipeOut(parsed_out_fifo);
   interface start = toPipeIn(start_fifo);
   interface done = toPipeOut(done_fifo);
endmodule

typedef enum {S0, S1, S2, S3} ParserState deriving (Bits, Eq);
instance FShow#(ParserState);
   function Fmt fshow (ParserState state);
      return $format(" State %x", state);
   endfunction
endinstance

(* synthesize *)
module mkParser(Parser);
   FIFOF#(EtherData) data_in_fifo <- mkSizedBypassFIFOF(4);
   FIFOF#(void) parse_done_fifo <- mkSizedFIFOF(1);

   ParseEthernet parse_ethernet <- mkParseEthernet();
   ParseIpv4 parse_ipv4 <- mkParseIpv4();

   mkConnection(parse_ethernet.unparsedOut, parse_ipv4.unparsedIn);

   let verbose = True;
   Reg#(Cycle_t) cycle <- mkReg(0);
   rule every;
      cycle <= cycle + 1;
   endrule

   Reg#(ParserState) curr_state <- mkReg(S0);

   // Parsing Graph
   (* fire_when_enabled *)
   rule state_S0 (curr_state == S0);
      let v = data_in_fifo.first;
      if (v.sop) begin
         curr_state <= S1;
         parse_ethernet.init;
         parse_ipv4.init;
         if (verbose) $display(fshow(cycle) + fshow("Done with") + fshow(curr_state));
      end
      else begin
         data_in_fifo.deq;
      end
   endrule
   (* fire_when_enabled *)
   rule state_S1 (curr_state == S1);
      let v <- toGet(parse_ethernet.done).get;
      curr_state <= S2;
      if (verbose) $display(fshow(cycle) + fshow("Done with") + fshow(curr_state));
   endrule
   (* fire_when_enabled *)
   rule state_S2 (curr_state == S2);
      let v <- toGet(parse_ipv4.done).get;
      curr_state <= S3;
      if (verbose) $display(fshow(cycle) + fshow("Done with") + fshow(curr_state));
   endrule
   (* fire_when_enabled *)
   rule state_S3 (curr_state == S3);
      let v <- toGet(data_in_fifo).get;
      if (verbose) $display(fshow(cycle) + fshow(curr_state));
      if (v.eop) begin
         curr_state <= S0;
         parse_ethernet.clear;
         parse_ipv4.clear;
         if (verbose) $display(fshow(cycle) + fshow("Done with") + fshow(curr_state));
      end
   endrule

   // Data dispatcher.
   rule state_S1_input (curr_state == S1);
      let v <- toGet(data_in_fifo).get;
      parse_ethernet.packetIn.enq(v.data);
      if (verbose) $display(fshow(cycle) + fshow("parse_ethernet enqueue ")+ fshow(v));
   endrule
   rule state_S2_input (curr_state == S2);
      let v <- toGet(data_in_fifo).get;
      parse_ipv4.packetIn.enq(v.data);
      if (verbose) $display(fshow(cycle) + fshow("parse_ipv4 enqueue ") + fshow(v));
   endrule

   // derive parse done from state machine
   interface frameIn = toPipeIn(data_in_fifo);
   interface parseDone = toPipeOut(parse_done_fifo);
endmodule

