// Copyright (c) 2016 Cornell University.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

typeclass StreamGearbox#(type ifc);
   
endtypeclass


instance StreamGearbox;
   module 
endinstance

// toHost

// toNetwork

// assume PacketDataT in host order
// m = 2n
function StreamerData#(m) combine(Vector#(2, StreamerData#(n)) v);
   StreamerData data = defaultValue;
   data.data = {v[1].data, v[0].data};
   data.mask = {v[1].mask, v[0].mask};
   data.sop = unpack(v[0].sop);
   data.eop = unpack(v[0].eop) || unpack(v[1].eop);
   return data;
endfunction

// rule handle sop

// rule handle odd flit

// rule handle even flit

