package Ethernet;

import EthMac                        ::*;
import EthPcs                        ::*;
import EthPma                        ::*;

instance Connectable#(MAC_XGMII, XGMII);


endinstance

endpackage
