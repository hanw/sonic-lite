// megafunction wizard: %LPM_MUX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_MUX 

// ============================================================
// File Name: xgmii_mux.v
// Megafunction Name(s):
// 			LPM_MUX
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module xgmii_mux (
	clock,
	data0x,
	data1x,
	data2x,
	data3x,
	sel,
	result);

	input	  clock;
	input	[65:0]  data0x;
	input	[65:0]  data1x;
	input	[65:0]  data2x;
	input	[65:0]  data3x;
	input	[1:0]  sel;
	output	[65:0]  result;

	wire [65:0] sub_wire0;
	wire [65:0] sub_wire5 = data3x[65:0];
	wire [65:0] sub_wire4 = data2x[65:0];
	wire [65:0] sub_wire3 = data1x[65:0];
	wire [65:0] result = sub_wire0[65:0];
	wire [65:0] sub_wire1 = data0x[65:0];
	wire [263:0] sub_wire2 = {sub_wire5, sub_wire4, sub_wire3, sub_wire1};

	lpm_mux	LPM_MUX_component (
				.clock (clock),
				.data (sub_wire2),
				.sel (sel),
				.result (sub_wire0)
				// synopsys translate_off
				,
				.aclr (),
				.clken ()
				// synopsys translate_on
				);
	defparam
		LPM_MUX_component.lpm_pipeline = 1,
		LPM_MUX_component.lpm_size = 4,
		LPM_MUX_component.lpm_type = "LPM_MUX",
		LPM_MUX_component.lpm_width = 66,
		LPM_MUX_component.lpm_widths = 2;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "1"
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "4"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "66"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "2"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: data0x 0 0 66 0 INPUT NODEFVAL "data0x[65..0]"
// Retrieval info: USED_PORT: data1x 0 0 66 0 INPUT NODEFVAL "data1x[65..0]"
// Retrieval info: USED_PORT: data2x 0 0 66 0 INPUT NODEFVAL "data2x[65..0]"
// Retrieval info: USED_PORT: data3x 0 0 66 0 INPUT NODEFVAL "data3x[65..0]"
// Retrieval info: USED_PORT: result 0 0 66 0 OUTPUT NODEFVAL "result[65..0]"
// Retrieval info: USED_PORT: sel 0 0 2 0 INPUT NODEFVAL "sel[1..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 66 0 data0x 0 0 66 0
// Retrieval info: CONNECT: @data 0 0 66 66 data1x 0 0 66 0
// Retrieval info: CONNECT: @data 0 0 66 132 data2x 0 0 66 0
// Retrieval info: CONNECT: @data 0 0 66 198 data3x 0 0 66 0
// Retrieval info: CONNECT: @sel 0 0 2 0 sel 0 0 2 0
// Retrieval info: CONNECT: result 0 0 66 0 @result 0 0 66 0
// Retrieval info: GEN_FILE: TYPE_NORMAL xgmii_mux.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL xgmii_mux.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL xgmii_mux.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL xgmii_mux.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL xgmii_mux_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL xgmii_mux_bb.v FALSE
// Retrieval info: LIB_FILE: lpm
