// altera_clkctrl.v

// Generated using ACDS version 14.0 200 at 2015.01.24.15:23:18

`timescale 1 ps / 1 ps
module altera_clkctrl (
		input  wire  inclk,  //  altclkctrl_input.inclk
		output wire  outclk  // altclkctrl_output.outclk
	);

	altera_clkctrl_altclkctrl_0 altclkctrl_0 (
		.inclk  (inclk),  //  altclkctrl_input.inclk
		.outclk (outclk)  // altclkctrl_output.outclk
	);

endmodule
