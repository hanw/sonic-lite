import PcieAlteraLIB ::*;


module mkPcieAlteraTestBench(Empty);


endmodule

